module handshake_p3(input clock, reset,
					input [3:0] ps2_data, input ps2_en,
					output [3:0] sound_code,	// Code for the music box
					input data_rq,		// Data request from music box
					output data_rd);		// Data ready for music box

// Your code goes here...

endmodule
