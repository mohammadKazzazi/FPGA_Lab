// 8-bit Adder/Subtractor datapath

module Part3(SW, LEDR, LEDG, KEY, HEX7, HEX6, HEX5, HEX4, HEX1, HEX0);
	input [8:0] SW;
	input [1:0] KEY;
	output [6:0] HEX7, HEX6, HEX5, HEX4, HEX1, HEX0;
	output [7:0] LEDR;
	output [8:0] LEDG;

	/* Your code goes here */
	
endmodule
