// Adder

module Part1(SW, LEDR, LEDG);
	input [8:0] SW;
	output [8:0] LEDR;
	output [4:0] LEDG;

	/* Your code goes here */

endmodule