`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/06/25 09:12:16
// Design Name: 
// Module Name: ram_read_write
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ram_read_write
    (
	 input              clk,
	 input              rst_n,
	 
     input      [31:0]  din,	 
	 output reg [31:0]  dout,
	 output reg         en,
	 output reg [3:0]   we,
	 output             rst,
	 output reg [31:0]  addr,
	 
	 input              start,
	 input      [31:0]  init_data,
	 output reg         start_clr,
	 output reg         write_end,
	 input      [31:0]  len,
	 input      [1:0]  freq
    );


assign rst = 1'b0 ;
	
localparam IDLE      = 3'd0 ;
localparam READ_RAM  = 3'd1 ;
localparam READ_END  = 3'd2 ;
localparam WRITE_RAM = 3'd3 ;
localparam WRITE_END = 3'd4 ;

reg [2:0] state ;
reg [9:0] len_tmp ;
reg [31:0] start_addr_tmp = 32'd0;
reg [15:0] sin_base [1023:0];
reg [9:0] read_ram_counter;

reg [9:0] write_ram_counter = 10'd1;


//write part	
always @(posedge clk or negedge rst_n)
begin
  if (~rst_n)
  begin
    state      <= IDLE  ;
	dout       <= 32'd0 ;
	en         <= 1'b0  ;
	we         <= 4'd0  ;
	addr       <= 32'd0 ;
	write_end  <= 1'b0  ;
	start_clr  <= 1'b0  ;
	len_tmp    <= 10'd0 ;
	start_addr_tmp <= 32'd0 ;
	read_ram_counter <= 10'd0;
	write_ram_counter <= 10'd1;
  end
	
  else
  begin
    case(state)
	IDLE            : begin
			            if (start)
						begin
			              state <= READ_RAM     ;
						  addr  <= 1'b0   ;
						  len_tmp <= len /(freq + 1) ;
						  dout <= init_data ;
						  en    <= 1'b1 ;
						  start_clr <= 1'b1 ;
						  read_ram_counter <= 10'd0;
						  write_ram_counter <= 10'd1;
						end			  
				        write_end <= 1'b0 ;
			          end

    
    READ_RAM        : begin
	                    if ((addr - start_addr_tmp) == len - 4)
						begin
						  state <= READ_END ;
						  en    <= 1'b0     ;
						end
						else
						begin
							sin_base[read_ram_counter] <= din; 
							read_ram_counter <= read_ram_counter + 1;
							addr <= addr + 32'd4;				

						end
						start_clr <= 1'b0 ;
					  end
					  
    READ_END        : begin
	                    addr  <= start_addr_tmp ;
	                    en <= 1'b1 ;
                        we <= 4'hf ;
					    state <= WRITE_RAM  ;					    
					  end
    
	WRITE_RAM       : begin
	                    if ((addr - start_addr_tmp) >= len_tmp - 4)
						begin
						  state <= WRITE_END ;
						  dout  <= 32'd0 ;
						  en    <= 1'b0  ;
						  we    <= 4'd0  ;
						end
						else
						begin
						  addr <= addr + 32'd4 ;
						  dout <= sin_base[write_ram_counter*(freq+1)] ;
						  write_ram_counter <= write_ram_counter+1;
						end
					  end
					  
	WRITE_END       : begin
	                    addr <= 32'd0 ;
						write_end <= 1'b1 ;
					    state <= IDLE ;					    
					  end	
	default         : state <= IDLE ;
	endcase
  end
end	
	
endmodule
