// BCD Counter

module Part4(CLOCK_50, KEY, HEX2, HEX1, HEX0);
	input CLOCK_50;
	input [0:0] KEY;
	output [6:0] HEX2, HEX1, HEX0;
	
	/* Your code goes here */
endmodule
